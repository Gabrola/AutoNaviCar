`ifndef _directions_vh_
`define _directions_vh_

`define None 3'd0
`define Forward 3'd1
`define Backward 3'd2
`define LForward 3'd3
`define RForward 3'd4
`define LBackward 3'd5
`define RBackward 3'd6

`endif